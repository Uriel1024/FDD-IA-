module gray ( 
	a,
	b,
	c,
	d,
	f,
	g,
	h,
	i
	) ;

input  a;
input  b;
input  c;
input  d;
inout  f;
inout  g;
inout  h;
inout  i;
