module sum_res ( 
	c1,
	op,
	a,
	b,
	s,
	cout,
	sel
	) ;

input  c1;
input  op;
input [3:0] a;
input [3:0] b;
inout [3:0] s;
inout  cout;
inout  sel;
