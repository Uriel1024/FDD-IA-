module sc ( 
	a,
	b,
	cin,
	sum,
	co
	) ;

input  a;
input  b;
input  cin;
inout  sum;
inout  co;
