module magnitud ( 
	a,
	b,
	c,
	d,
	f,
	g,
	h
	) ;

input  a;
input  b;
input  c;
input  d;
inout  f;
inout  g;
inout  h;
