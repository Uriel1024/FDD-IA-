module dec ( 
	e,
	d
	) ;

input [3:0] e;
inout [9:0] d;
