module cod ( 
	e,
	s,
	con,
	y
	) ;

input [8:0] e;
inout [2:0] s;
input  con;
inout  y;
