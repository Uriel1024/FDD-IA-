module dec ( 
	e,
	d
	) ;

input [4:0] e;
inout [9:0] d;
