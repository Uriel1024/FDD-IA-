module mux_8a1 ( 
	i0,
	i1,
	i2,
	i3,
	i4,
	i5,
	i6,
	i7,
	s,
	y
	) ;

input  i0;
input  i1;
input  i2;
input  i3;
input  i4;
input  i5;
input  i6;
input  i7;
input [2:0] s;
inout  y;
