module p11_mux ( 
	a,
	b,
	c,
	d,
	x,
	y,
	z,
	f
	) ;

input  a;
input  b;
input  c;
input  d;
input  x;
input  y;
input  z;
inout  f;
