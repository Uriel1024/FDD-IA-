module m_sum ( 
	a,
	b,
	sum,
	cout
	) ;

input  a;
input  b;
inout  sum;
inout  cout;
