module display ( 
	a,
	b,
	c,
	d,
	f,
	g,
	h,
	i,
	j,
	k,
	l
	) ;

input  a;
input  b;
input  c;
input  d;
inout  f;
inout  g;
inout  h;
inout  i;
inout  j;
inout  k;
inout  l;
