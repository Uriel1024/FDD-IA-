module display ( 
	e,
	dis
	) ;

input [4:0] e;
inout [6:0] dis;
