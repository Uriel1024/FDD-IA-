module bcd ( 
	e,
	dis
	) ;

input [3:0] e;
inout [6:0] dis;
