module sumadordosbits ( 
	a,
	b,
	cin,
	sum,
	cout
	) ;

input [1:0] a;
input [1:0] b;
input  cin;
inout [1:0] sum;
inout  cout;
