module resta ( 
	a,
	b,
	pi,
	resta,
	po
	) ;

input  a;
input  b;
input  pi;
inout  resta;
inout  po;
