module cod ( 
	e,
	s,
	y
	) ;

input [7:0] e;
inout [2:0] s;
inout  y;
